LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FFD IS
PORT (
		ENT: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		CLK,RST,ENABLE: IN STD_LOGIC;
		SD:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END FFD;

ARCHITECTURE FFD_ARCH OF FFD IS
BEGIN
	PROCESS(CLK,RST)
	BEGIN
		IF RST ='1' THEN
			SD <="00000000";
		ELSIF CLK'EVENT AND CLK='1' THEN
			IF ENABLE ='1' THEN
				SD <= ENT;
			END IF;
		END IF;
	END PROCESS;
END FFD_ARCH;
