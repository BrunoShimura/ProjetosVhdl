LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY pand IS
	PORT(
		E1: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		E2: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		S: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
	
END pand;

ARCHITECTURE pand_arch OF pand IS

BEGIN
	S <= E1 + E2;
END pand_arch ;
